module i5SEXT (
input [5:0] s_in,
output [15:0] s_out
);

endmodule

// QUICK AND DIRTY: ONLY WORKS UP TO 4-INPUT MUX
module o16MUX21 
(input Sel;
input [15:0] i_data [X];
output [15:0] o_data;
);

case(Sel)
	
endmodule

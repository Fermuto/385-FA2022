module CPU (
);
endmodule

module Status (
);

endmodule

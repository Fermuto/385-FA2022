module compute 
endmodule

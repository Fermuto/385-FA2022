module Instruction {
);

endmodule

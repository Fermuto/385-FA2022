module IR (
);
endmodule

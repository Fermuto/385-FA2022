
module lab61soc (
	clk_clk);	

	input		clk_clk;
endmodule

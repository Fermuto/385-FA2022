module ALU (
);

endmodule
module MDR (
);
endmodule
module i11SEXT (
input [10:0] s_in,
output [15:0] s_out
);

endmodule
module multiplier (input logic Clk, Reset_Load_Clear, Run, 
				input logic [7:0] SW,
				output logic [7:0] Aval, Bval,
				output logic Xval,
				output logic [6:0] HEX0, 
										 HEX1, 
										 HEX2, 
										 HEX3, 
										 HEX4,
										 HEX5

);

endmodule

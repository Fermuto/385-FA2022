module i9SEXT (
input [8:0] s_in,
output [15:0] s_out
);

endmodule
module MAR (
);

endmodule
/************************************************************************
Avalon-MM Interface VGA Text mode display

Register Map:
0x000-0x0257 : VRAM, 80x30 (2400 byte, 600 word) raster order (first column then row)
0x258        : control register

VRAM Format:
X->
[ 31  30-24][ 23  22-16][ 15  14-8 ][ 7    6-0 ]
[IV3][CODE3][IV2][CODE2][IV1][CODE1][IV0][CODE0]

IVn = Draw inverse glyph
CODEn = Glyph code from IBM codepage 437

Control Register Format:
[[31-25][24-21][20-17][16-13][ 12-9][ 8-5 ][ 4-1 ][   0    ] 
[[RSVD ][FGD_R][FGD_G][FGD_B][BKG_R][BKG_G][BKG_B][RESERVED]

VSYNC signal = bit which flips on every Vsync (time for new frame), used to synchronize software
BKG_R/G/B = Background color, flipped with foreground when IVn bit is set
FGD_R/G/B = Foreground color, flipped with background when Inv bit is set

************************************************************************/
`define NUM_REGS 601 //80*30 characters / 4 characters per register
`define CTRL_REG 600 //index of control register

module vga_text_avl_interface (
	// Avalon Clock Input, note this clock is also used for VGA, so this must be 50Mhz
	// We can put a clock divider here in the future to make this IP more generalizable
	input logic CLK,
	
	// Avalon Reset Input
	input logic RESET,
	
	// Avalon-MM Slave Signals
	input  logic AVL_READ,					// Avalon-MM Read
	input  logic AVL_WRITE,					// Avalon-MM Write
	input  logic AVL_CS,					// Avalon-MM Chip Select
	input  logic [3:0] AVL_BYTE_EN,			// Avalon-MM Byte Enable
	input  logic [9:0] AVL_ADDR,			// Avalon-MM Address
	input  logic [31:0] AVL_WRITEDATA,		// Avalon-MM Write Data
	output logic [31:0] AVL_READDATA,		// Avalon-MM Read Data
	
	// Exported Conduit (mapped to VGA port - make sure you export in Platform Designer)
	output logic [3:0]  red, green, blue,	// VGA color channels (mapped to output pins in top-level)
	output logic hs, vs						// VGA HS/VS
);

logic [31:0] LOCAL_REG       [601]; // Registers
//put other local variables here
logic vssig, blank, sync, VGA_Clk;
logic [9:0] drawxsig, drawysig, spritexsig, spriteysig;
logic [9:0] c_div, r_div, f_addr, reg_base;
logic [1:0] reg_sp;
logic [31:0] grab_reg;
logic [7:0] char_code;
logic [3:0] Fore_R, Fore_B, Fore_G, Back_R, Back_B, Back_G;

logic [10:0] sprite_addr;
logic [7:0] sprite_data, sprite_out;
//Declare submodules..e.g. VGA controller, ROMS, etc

	
vga_controller controller0(.Clk (CLK), .Reset (RESET), .hs (hs), .vs (vs), .pixel_clk (VGA_Clk), .blank (blank), .sync (sync), .DrawX (drawxsig), .DrawY (drawysig));

font_rom bitmaps (.addr (sprite_addr), .data (sprite_out));

   
// Read and write from AVL interface to register block, note that READ waitstate = 1, so this should be in always_ff
always_ff @(posedge CLK) begin
	if (AVL_CS && AVL_READ)
	begin
		AVL_READDATA <= LOCAL_REG[AVL_ADDR];
	end
	
	else if (AVL_CS && AVL_WRITE)
	begin
		case (AVL_BYTE_EN)
		4'b1111:
			begin
				LOCAL_REG[AVL_ADDR] <= AVL_WRITEDATA;
			end
		4'b1100:
			begin
				LOCAL_REG[AVL_ADDR][31:16] <= AVL_WRITEDATA[31:16];
			end
		4'b0011:
			begin
				LOCAL_REG[AVL_ADDR][15:0] <= AVL_WRITEDATA[15:0];
			end
		4'b1000:
			begin
				LOCAL_REG[AVL_ADDR][31:24] <= AVL_WRITEDATA[31:24];
			end
		4'b0100:
			begin
				LOCAL_REG[AVL_ADDR][23:16] <= AVL_WRITEDATA[23:16];
			end
		4'b0010:
			begin
				LOCAL_REG[AVL_ADDR][15:8] <= AVL_WRITEDATA[15:8];
			end
		4'b0001:
			begin
				LOCAL_REG[AVL_ADDR][7:0] <= AVL_WRITEDATA[7:0];
			end
		endcase
	end
end


//handle drawing (may either be combinational or sequential - or both).

always_ff @(VGA_Clk)
begin
	if (blank == 1'b0)
	begin
		red <= 4'h0;
		green <= 4'h0;
		blue <= 4'h0;
	end
	
	else
	begin
		c_div <= (drawxsig >> 3); // divide by 8
		r_div <= (drawxsig >> 4); // divide by 16

		f_addr <= (r_div * 8'd80) + c_div; //flatten 2d coords to 1d
		
		reg_base <= (f_addr >> 2);
		reg_sp <= (f_addr % 4);
		
		grab_reg <= LOCAL_REG[reg_base]; //grab character hex code
		case (reg_sp)
		2'b00:char_code <= grab_reg[7:0];
		2'b01:char_code <= grab_reg[15:8];
		2'b10:char_code <= grab_reg[23:16];
		2'b11:char_code <= grab_reg[31:24];
		endcase
		
		spritexsig <= (c_div * 8'd8); // determine top left corner of sprite
		spriteysig <= (r_div * 8'd16);
		
		sprite_addr = (drawysig - spriteysig + (16 * char_code));
		
		Fore_R <= LOCAL_REG[600][24:21];
		Fore_G <= LOCAL_REG[600][20:17];
		Fore_B <= LOCAL_REG[600][16:13];
		Back_R <= LOCAL_REG[600][12:9];
		Back_G <= LOCAL_REG[600][8:5];
		Back_B <= LOCAL_REG[600][4:1];
		
		for (int i = 0; i < $size(sprite_out); i++)
			sprite_data[7-i] <= sprite_out[i];
		
		if (sprite_data[drawxsig - spritexsig] == 1'b1)
		begin
			red = Fore_R;
			green = Fore_G;
			blue = Fore_B;
		end
		
		else
		begin
			red = Back_R;
			green = Back_G;
			blue = Back_B;
		end
	end
	
end

endmodule
